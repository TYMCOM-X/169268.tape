ARLINGTON  5632 1590
ATLANTA    7260 2083
BALTIMORE  5510 1575
BIRMINGHAM 7518 2446
BOISE      7096 7869
BOSTON     4422 1249
BUFFALO    5075 2326
CARSONCITY 8139 8306
CHICAGO    5986 3426
COLUMBUS   5972 2555
CUPERTINO  8583 8619
DALLAS     8436 4034
DENVER     7501 5899
DESMOINES  6471 4275
DETROIT    5536 2828
DURHAM     6331 1499
HARTFORD   4687 1373
HOUSTON    8938 3536
LOSANGELES 9213 7878
LOUISVILLE 6529 2772
LYNDHURST  4993 1433
MEMPHIS    7471 3125
MIAMI      8351  527
MILWAUKEE  5788 3589
MINNEAPOLS 5777 4513
NEWORLEANS 8483 2638
NEWYORK    4997 1406
OKLACITY   7947 4373
OMAHA      6687 4595
PHILA      5251 1458
PHOENIX    9135 6748
PORTLAND   6799 8914
ROCHESTER  4913 2195
SALTLAKE   7576 7065
SANFRAN    8492 8719
SEATTLE    6336 8896
STLOUIS    6807 3482
SYRACUSE   4798 1990
VALLEYFRG  5250 1515
WICHITA    7489 4520
