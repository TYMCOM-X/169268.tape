From Mallek Khellaf (922-7089)
To   Rick Della Rocco


Present 56 kb links in TYMNET
=====================================================
City1           ST NPA NXX City2           ST NPA NXX
=====================================================
NORRISTOWN      PA 215 666 NEWARK          NJ 201 824 
NORRISTOWN      PA 215 666 FAIRFAX         VA 703 691 
NORRISTOWN      PA 215 666 SAN JOSE        CA 408 433 
NORRISTOWN      PA 215 666 HAZELWOOD       MO 314 232 
NORRISTOWN      PA 215 666 DALLAS          TX 214 637 
DALLAS          TX 214 637 SAN FRANCISCO   CA 415 896 
DALLAS          TX 214 637 SAN JOSE        CA 408 433 
DALLAS          TX 214 637 SAN JOSE        CA 408 433 
DALLAS          TX 214 637 MINNEAPOLIS     MN 612 333 
DALLAS          TX 214 637 NEWARK          NJ 201 824 
FREMONT         CA 415 498 DALLAS          TX 214 637 
FREMONT         CA 415 498 FREMONT         CA 415 498 
FREMONT         CA 415 498 FREMONT         CA 415 498 
FREMONT         CA 415 498 FREMONT         CA 415 498 
FREMONT         CA 415 498 FREMONT         CA 415 498 
FREMONT         CA 415 498 FREMONT         CA 415 498 
FREMONT         CA 415 498 FREMONT         CA 415 498 
FREMONT         CA 415 498 CHICAGO         IL 312 427 
FREMONT         CA 415 498 SAN FRANCISCO   CA 415 543 
FREMONT         CA 415 498 SAN JOSE        CA 408 433 
FREMONT         CA 415 498 SAN JOSE        CA 408 433 
FREMONT         CA 415 498 SAN JOSE        CA 408 433 
FREMONT         CA 415 498 VERNON          CA 213 589 
NEWARK          NJ 201 824 FAIRFAX         VA 703 691 
NEWARK          NJ 201 824 CHICAGO         IL 312 427 
NEWARK          NJ 201 824 BOSTON          MA 617 439 
NEWARK          NJ 201 824 DORAVILLE       GA 404 451 
SAN FRANCISCO   CA 415 896 HONOLULU        HI 808 531 
SAN FRANCISCO   CA 415 896 HONOLULU        HI 808 531 
DENVER          CO 303 860 DALLAS          TX 214 637 
BALTIMORE       MD 301 685 FAIRFAX         VA 703 691 
FAIRFAX         VA 703 691 DALLAS          TX 214 637 
FAIRFAX         VA 703 691 ROCKVILLE       MD 301 840 
FAIRFAX         VA 703 691 SAN FRANCISCO   CA 415 543 
FAIRFAX         VA 703 691 HOUSTON         TX 713 497 
FAIRFAX         VA 703 691 DORAVILLE       GA 404 451 
SEATTLE         WA 206 284 SAN FRANCISCO   CA 415 543 
NEWPORT BEACH   CA 714 756 SAN DIEGO       CA 619 560 
NEWPORT BEACH   CA 714 756 SAN FRANCISCO   CA 415 896 
NEWPORT BEACH   CA 714 756 SAN JOSE        CA 408 433 
NEWPORT BEACH   CA 714 756 VERNON          CA 213 589 
NEWPORT BEACH   CA 714 756 NEWARK          NJ 201 824 
NEWPORT BEACH   CA 714 756 DALLAS          TX 214 637 
CHICAGO         IL 312 427 DENVER          CO 303 860 
CHICAGO         IL 312 427 FAIRFAX         VA 703 691 
CHICAGO         IL 312 427 BOSTON          MA 617 439 
CHICAGO         IL 312 427 SAN FRANCISCO   CA 415 543 
CHICAGO         IL 312 427 SAN JOSE        CA 408 433 
CHICAGO         IL 312 427 SAN JOSE        CA 408 433 
CHICAGO         IL 312 427 MINNEAPOLIS     MN 612 333 
CHICAGO         IL 312 427 PLYMOUTH        MI 313 455 
CHICAGO         IL 312 427 DETROIT         MI 313 963 
CHICAGO         IL 312 427 DALLAS          TX 214 637 
CHICAGO         IL 312 427 DALLAS          TX 214 637 
BOSTON          MA 617 439 FAIRFAX         VA 703 691 
SAN FRANCISCO   CA 415 543 SAN JOSE        CA 408 433 
SAN JOSE        CA 408 433 NEWARK          NJ 201 824 
SAN JOSE        CA 408 433 DALLAS          TX 214 637 
MISSION         KS 913 384 DALLAS          TX 214 637 
PLYMOUTH        MI 313 455 FAIRFAX         VA 703 691 
PLYMOUTH        MI 313 455 DETROIT         MI 313 963 
HAZELWOOD       MO 314 232 FAIRFAX         VA 703 691 
HAZELWOOD       MO 314 232 CHICAGO         IL 312 427 
HAZELWOOD       MO 314 232 DALLAS          TX 214 637 
VERNON          CA 213 589 DALLAS          TX 214 637 
HOUSTON         TX 713 497 DALLAS          TX 214 637 
DALLAS          TX 214 637 MIAMI           FL 305 477 
DORAVILLE       GA 404 451 DALLAS          TX 214 637 
  