ALBANY         4639 1629
ALBUQUERQU     8549 5887
ALEXANDRIA     8409 3168
ALLEN PARK     5536 2828
ALTOONA        5460 1972
AMARILLO       8266 5076
ANN ARBOR      5602 2918
ASHEVILLE      6749 2001
ASPINWALL      5621 2185
ATLANTA        7260 2083
AUGUSTA        7089 1674
AUSTIN         9005 3996
BALTIMORE      5510 1575
BATAVIA        4993 2250
BATH           5033 2052
BATTLE CRE     5713 3124
BAY PINES      8224 1159
BECKLEY        6218 2043
BEDFORD        4424 1283
BIG SPRING     8847 4800
BILOXI         8296 2481
BIRMINGHAM     7518 2446
BOISE          7096 7869
BONHAM         8234 3996
BOSTON         4431 1254
BRAINTREE      4440 1222
BRECKSVILL     5604 2515
BROCKTON       4465 1205
BRONX          4997 1406
BROOKLYN       4997 1406
BUFFALO        5075 2326
BUTLER         5534 2221
CANANDAIGU     4931 2117
CASTLE POI     4861 1504
CHARLESTON     7021 1281
CHEYENNE       7203 5958
CHICAGO        5986 3426
CHILLICOTH     6088 2480
CINCINNATI     6263 2679
CLARKSBURG     5865 2095
CLEVELAND      5574 2543
COATESVILL     5310 1553
COLUMBIA       6901 1589
COLUMBUS       5972 2555
DALLAS         8436 4034
DANVILLE       6322 3245
DAYTON         6113 2705
DECATUR        7260 2083
DENVER         7501 5899
DES MOINES     6471 4275
DETROIT        5536 2828
DUBLIN         7354 1718
DURHAM         6331 1499
EAST ORANG     5015 1442
EL PASO        9231 5655
ERIE           5321 2397
FARGO          5615 5182
FAYETTEVIL     7600 3872
FORT WAYNE     5942 2982
FRESNO         8669 8239
FT HARRISO     6336 7348
FT HOWARD      5513 1548
FT LYON        7756 5501
FT MEADE       6463 5966
FT. HARRIS     6336 7348
GAINESVILL     7838 1310
GRAND ISLA     6901 4936
GRAND JUNC     7804 6438
GRAND PRAR     8458 4066
HAMPTON        5891 1252
HARTFORD       4687 1373
HINES          6001 3455
HOT SPRING     6666 5898
HOUSTON        8938 3536
HUNTINGTON     6212 2299
INDIANAPOL     6272 2992
IOWA CITY      6313 3972
IRON MOUNT     5266 3890
JACKSON        8035 2880
KANSAS CIT     7027 4203
KERRVILLE      9143 4226
KNOXVILLE      6490 4172
LAKE CITY      7768 1419
LAKEWOOD       7507 5912
LAS VEGAS      8665 7411
LEAVENWORT     7008 4272
LEBANON        5304 1679
LEXINGTON      6459 2562
LINCOLN        6823 4674
LITTLE ROC     7721 3451
LIVERMORE      8504 8606
LOMA LINDA     9183 7711
LONG BEACH     9271 7856
LOS ANGELE     9218 7914
LOUISVILLE     6529 2772
LYONS          5061 1468
MADISON        5887 3796
MANCHESTER     4354 1388
MARION         6882 3202
MARLIN         8739 3931
MARTINEZ       8438 8677
MARTINSBUR     5611 1783
MEMPHIS        7471 3125
MIAMI          8351  527
MILES CITY     6155 6433
MINNEAPOLI     5777 4513
MONTEREY       8743 8601
MONTGOMERY     7692 2247
MONTROSE       4894 1470
MOUNTAIN H     6594 2051
MURFREESBO     7036 2618
MUSKOGEE       7746 4042
N. LITTLE      7721 3451
NASHVILLE      7010 2710
NEW ORLEAN     8483 2638
NEW YORK       4997 1406
NEWARK         5015 1430
NEWINGTON      4705 1368
NORTH CHIC     5909 3503
NORTHAMPTO     4587 1442
NORTHPORT      4904 1342
OKLAHOMA C     7947 4373
OMAHA          6687 4595
PALO ALTO      8562 8668
PERRY POIN     5411 1533
PHILADELPH     5251 1458
PHOENIX        8983 7203
PITTSBURGH     5621 2185
POPLAR BLU     7184 3333
PORTLAND       6799 8914
PRESCOTT       8917 6872
PROVIDENCE     4550 1219
RENO           8064 8323
RICHMOND       5906 1472
ROANOKE        6196 1801
ROMNEY         5706 1878
ROSEBURG       7318 8982
SAGINAW        5404 3074
SALEM          6196 1801
SALISBURY      6540 1691
SALT LAKE      7576 7065
SAN ANTONI     9209 4088
SAN DIEGO      9445 7657
SAN FRANCI     8492 8719
SEATTLE        6336 8896
SEPULVEDA      9168 7922
SHERIDAN       6535 6505
SHREVEPORT     8272 3495
SIOUX FALL     6279 4900
SPOKANE        6247 8180
ST. CLOUD      5721 4705
ST. LOUIS      6842 3492
ST. PAUL       5777 4513
ST. PETERS     8224 1159
SYRACUSE       4798 1990
TACOMA         6415 8906
TAMPA          8173 1147
TEMPLE         8812 3992
TOGUS          3961 1370
TOMAH          5792 4042
TOPEKA         7110 4369
TROY           4639 1629
TUCSON         9345 6485
TUSCALOOSA     7643 2535
TUSKEGEE       7628 2153
W. LOS ANG     9218 7914
WACO           8706 3993
WALLA WALL     6611 8269
WASHINGTON     5622 1583
WEST HAVEN     4800 1340
WHITE CITY     7480 8889
WHITE RIVE     4327 1585
WICHITA        7489 4520
WILKES-BAR     5093 1723
WILMINGTON     5326 1485
WINSTON-SA     6440 1710
    