
(ENFE:33,39)NEWFAX.CKT                                       TABS 9,29,41,50,57


                    TELCO  CIRCUIT  INSTALLATION  LOG
                    ---------------------------------
                                                         TERMINATION  POINT
LINE    CIRCUIT NUMBER      DATE INST.  VENDOR   TECH       AND/OR REQ #
===============================================================================
   1 |  36 LGGS 61323     | 02/28/84  | C & P  | KRJ  | C 0781477
-------------------------------------------------------------------------------
   2 |  36 LGGS 61470     | 02/29/84  | C & P  | CG   | C 078435
-------------------------------------------------------------------------------
   3 |  36 FDDA 25671     | 03/27/84  | C & P  | CG   | N 2891969  2WR FTCC
-------------------------------------------------------------------------------
   4 |  36 FDDA 25756     | 03/27/84  | C & P  | CG   | "    "    "    "
-------------------------------------------------------------------------------
   5 |  36 FDDA 25757     | 03/27/84  | C & P  | CG   | "    "    "    "
-------------------------------------------------------------------------------
   6 |  36 LGFS 77271     | 03/28/84  | C & P  | TD   | C 0875978
-------------------------------------------------------------------------------
   7 |  36 LFGS 69590     | 03/29/84  | C & P  | TD   | C 0876584
-------------------------------------------------------------------------------
   8 |  36 LGGS 68271     | 03/29/84  | C & P  | TD   | C 0785531
-------------------------------------------------------------------------------
   9 |  36 LGGS 77291     | 03/29/84  | C & P  | TD   | C 0875999
-------------------------------------------------------------------------------
  10 |  352-8885          | 04/02/84  | C & P  | BF   | N 2891959
-------------------------------------------------------------------------------
  11 |  352-8886          | 04/02/84  | C & P  | BF   | "    "    "    "
-------------------------------------------------------------------------------
  12 |  352-8887          | 04/02/84  | C & P  | BF   | "    "    "    "
-------------------------------------------------------------------------------
  13 |  36 LGFS 77269     | 04/02/84  | C & P  | JT   | C 0875976
-------------------------------------------------------------------------------
  14 |  36 LGGS 77273     | 04/03/84  | C & P  | KRJ  | C 0875980
-------------------------------------------------------------------------------
  15 |  36 LGFS 77275     | 04/04/84  | C & P  | KRJ  | C 0875982
-------------------------------------------------------------------------------
  16 |  36 LGGS 69069     | 04/16/84  | C & P  | FH   | C 0797488
-------------------------------------------------------------------------------
  17 |  36 FDDA 27820     | 04/16/84  | C & P  | GGS  | N 2892556
-------------------------------------------------------------------------------
  18 |  36 FDDA 27821     | 04/17/84  | C & P  | KRJ  | N 2892557 19;5
-------------------------------------------------------------------------------
  19 |  36 FDEA 27759     | 04/20/84  | C & P  | FLH  | C 2903154 2WR 22;7
-------------------------------------------------------------------------------
  20 |  36 LGGS 77292     | 04/26/84  | C & P  | KRJ  | FDEA 608117   25;8
-------------------------------------------------------------------------------
  21 |  36 LGFS 70210     | 04/30/84  | C & P  | CHUCK| FDEA 552666   25;9
-------------------------------------------------------------------------------
  22 |  FDEA 503333       | 05/02/84  | C & P  |TOM D.| C 0884036     25;10
-------------------------------------------------------------------------------
  23 |  FDEA 552665       | 05/02/84  | C & P  |TOM D.| C 0888053     25;11
-------------------------------------------------------------------------------
  24 |  36 LGGS 60910     | 05/10/84  | C & P  | CG   | FDEA 713854   21;4
-------------------------------------------------------------------------------
  25 |  36 LGFS 64442     | 05/14/84  | C & P  | KRJ  | FDEA 724027   25;12
-------------------------------------------------------------------------------
  26 |  36 LGGS 15733     | 05/25/84  | C & P  | CG   | FDEA 552710   MV'D-22;2
-------------------------------------------------------------------------------











-------------------------------------------------------------------------------
  27 |  36 LGFS 70908     | 06/12/84  | C & P  | CG   | FDEA 50331     4;6
-------------------------------------------------------------------------------
  28 |  36 FDEA 28099     | 06/14/84  | C & P  | CG   | C2904296  2WR 22;8
-------------------------------------------------------------------------------
  29 |  36 FDEA 28555     | 06/27/84  | C & P  | CG   | N2908978       2;4
-------------------------------------------------------------------------------
  30 |  36 FD   28532     | 06/--/84  | C & P  |      |                2;3
-------------------------------------------------------------------------------
  31 |  36 LGGS 66894 CD  | 06/29/84  | C & P  | NH   | FDEA 363546    2;6
-------------------------------------------------------------------------------
  32 |  36 FDDA 28607     | 07/02/84  | C & P  | CG   | N3397660       2;7
-------------------------------------------------------------------------------
  33 |  36 FDEA 28613     | 07/02/84  | C & P  | CG   | N3398129  2WR 22;9
-------------------------------------------------------------------------------
  34 |  36 LGGS 66892     | 07/03/84  | C & P  | CG   | FDEA 362951    2;5
-------------------------------------------------------------------------------
  35 |  691-0036 & 0037   | 07/03/84  | C & P  | VAF  | STAND ALONE DATA JACKS
-------------------------------------------------------------------------------
  36 |  36 LGFS 67018     | 07/05/84  | C & P  | FH   | C0892062      25;1
-------------------------------------------------------------------------------
  37 |  36 LGFS 65347     | 07/11/84  | C & P  | FH   | FDEA 358081  25;6
-------------------------------------------------------------------------------
  38 |  36 LGFS 67686     | 07/12/84  | C & P  | CG   | FDEA 367213  25;4
-------------------------------------------------------------------------------
  39 |  36 LGFS 79761     | 07/12/84  | C & P  | CG   | FDEA 364540  25;5
-------------------------------------------------------------------------------
  40 |  36 LGFS 67694     | 07/17/84  | C & P  | CG   | FDEA 368367  2;8
-------------------------------------------------------------------------------
  41 |  36 FDDA 28876     | 07/20/84  | C & P  | CG   | N3400082     3;1
-------------------------------------------------------------------------------
  42 |  36 FDEA 28613     | 08/10/84  | C & P  | FH   | N3398129     22;9
-------------------------------------------------------------------------------
  43 |  36 FDEA 28714     | 08/15/84  | C & P  | PHIL | N3398139     26;2
-------------------------------------------------------------------------------
  44 |  36 FDEA 28715     | 08/15/84  | C & P  | PHIL | N3398140     26;3
-------------------------------------------------------------------------------
  45 |  36 FDEA 28716     | 08/15/84  | C & P  | PHIL | N3398141     26;4
-------------------------------------------------------------------------------
  46 |  36 FDEA 28717     | 08/15/84  | C & P  | PHIL | N3398142     26;5
-------------------------------------------------------------------------------
  47 |  36 FDEA 29161     | 08/16/84  | C & P  | MTW  | N3764445      3;3
-------------------------------------------------------------------------------
  48 |  36 LGFS 80574     | 08/21/84  | C & P  | KRJ  | FDEA 372775  26;6
-------------------------------------------------------------------------------
  49 |  36 FDEA 28718     | 08/21/84  | C & P  | KRJ  | N3398143     26;7
-------------------------------------------------------------------------------
  50 |  36 FDEA 28719     | 08/22/84  | C & P  | KRJ  | N3398144     26;8
-------------------------------------------------------------------------------
  51 |  36 FDEA 29285     | 08/28/84  | C & P  | KRJ  | N3764492      3;2
-------------------------------------------------------------------------------
  52 |  36 FDEA 29110     | 08/29/84  | C & P  | KRJ  | N2925820      3;4
-------------------------------------------------------------------------------
  53 |  36 LGGS 80467     | 08/29/84  | C & P  | KRJ  | FDEA 372774  26;10
-------------------------------------------------------------------------------









-------------------------------------------------------------------------------
  54 |  36 LGGS 80438     | 08/29/84  | C & P  | KRJ  | FDEA 695766  26;9
-------------------------------------------------------------------------------
  55 |  36 FDDA 29304     | 08/29/84  | C & P  | KRJ  | N3775478     13;2
-------------------------------------------------------------------------------
  56 |  36 XGGS 81820     | 08/31/84  | C & P  | CMG  | DIALNET RJ21;5 & 6
-------------------------------------------------------------------------------
  57 |  36 XGGS 81806     | 08/31/84  | C & P  | CMG  | DIALNET RJ21;3 & 4
-------------------------------------------------------------------------------
  58 |  36 LGFS 66624     | 09/05/84  | C & P  | KRJ  | FDEA 367215   3;8
-------------------------------------------------------------------------------
  59 |  36 LGFS 66285     | 09/05/84  | C & P  | KRJ  | FDES 361779.001 22;10
-------------------------------------------------------------------------------
  60 |  36 LGFS 80579     | 09/12/84  | C & P  | KRJ  | FDEA 695767  26;1
-------------------------------------------------------------------------------
  61 |  36 XGGS 8192/DDS  | 09/12/84  | C & P  | KRJ  | C 0945935    DDS CAB.
-------------------------------------------------------------------------------
  62 |  36 LGFS 82033     | 09/13/84  | C & P  | KRJ  | FDEA 220964  SLOT 1
-------------------------------------------------------------------------------
  63 |  36 FDEA 29416     | 09/13/84  | C & P  | KRJ  | N 3764499    SLOT 2
-------------------------------------------------------------------------------
  64 |  36 FDEA 29446     | 09/13/84  | C & P  | KRJ  | N 3764508    SLOT 3
-------------------------------------------------------------------------------
  65 |  36 LGGS 81458     | 09/13/84  | C & P  | KRJ  | FDEC 002812.013 SLOT 4
-------------------------------------------------------------------------------
  66 |  36 LGFS 81548     | 09/13/84  | C & P  | KRJ  | FDEA 899712  SLOT 5
-------------------------------------------------------------------------------
  67 |  36 LGGS 80611     | 09/13/84  | C & P  | KRJ  | FDEA 372776  SLOT 6
-------------------------------------------------------------------------------
  68 |  36 FDDA 29197     | 09/17/84  | C & P  | KRJ  | N 3399865    SLOT 7
-------------------------------------------------------------------------------
  69 |  36 FDDA 29198     | 09/17/84  | C & P  | KRJ  | N 3399866    SLOT 8
-------------------------------------------------------------------------------
  70 |  36 FDDA 29196     | 09/17/84  | C & P  | KRJ  | N 3399870B   SLOT 9
-------------------------------------------------------------------------------
  71 |  36 FDDA 29507     | 09/24/84  | C & P  | KRJ  | N 3765915    SLOT 10
-------------------------------------------------------------------------------
  72 |  36 LGFS 80954     | 09/26/84  | C & P  | KRJ  | FDEA 374279  SLOT 11
-------------------------------------------------------------------------------
  73 |  36 FDEA 29547     | 09/27/84  | C & P  | KRJ  | C 3765420    SLOT 12
-------------------------------------------------------------------------------
  74 |  36 FDEA 29067     | 10/03/84  | C & P  | KRJ  | N 3398170    SLOT 12
-------------------------------------------------------------------------------
  75 |  36 LGFS 84373     | 10/10/84  | C & P  | KRJ  | FDEA 380172  SLOT 13
-------------------------------------------------------------------------------
  76 |  36 LGFS 84511     | 10/10/84  | C & P  | KRJ  | FDEA 380173  SLOT 14
-------------------------------------------------------------------------------
  77 |  36 FDEA 29713CD   | 10/25/84  | C & P  | HJPO | N 3767187    SLOT 15
-------------------------------------------------------------------------------
  78 |  36 FDDA 29698     | 10/29/84  | C & P  | KRJ  | C 3765446      23;1
-------------------------------------------------------------------------------
  79 |  36 FDDA 29842     | 11/09/84  | C & P  | HJPO | N 3767360    SLOT 16
-------------------------------------------------------------------------------
  80 |  36 LGGC 150378    | 11/14/84  | C & P  | KRJ  | N 3767228    SLOT 17
-------------------------------------------------------------------------------
  81 |  36 LGGC 150379    | 11/15/84  | C & P  | KRJ  | N 3767230    SLOT 18
-------------------------------------------------------------------------------
  82 |  36 LGGS 105384    | 11/19/84  | C & P  | GGS  | N 3767375    SLOT 19
-------------------------------------------------------------------------------








-------------------------------------------------------------------------------
  83 |  36 FDEA 29534 CD  | 11/19/84  | C & P  | GGS  | C 3765417 B CANCELLED
-------------------------------------------------------------------------------
  84 |  36 LGGS 150385    | 11/19/84  | C & P  | GGS  | N 3767384    SLOT 21
-------------------------------------------------------------------------------
  85 |  36 LGGC 151854    | 11/30/84  | C & P  | KRJ  | N 3765533    SLOT 22
-------------------------------------------------------------------------------
  86 |  36 FDDA 28876     | 12/14/84  | C & P  | CG   | D3770393 DISC @3 SLOT1
-------------------------------------------------------------------------------
  87 |  301-293-1201      | 12/17/84  | C & P  | MTW  | C 0965127 BLOK BK WALL
-------------------------------------------------------------------------------
  88 |  36 XGGS 89957     | 12/19/84  | C & P  | TD   | C 0963151  DIGITAL CAB.
-------------------------------------------------------------------------------
  89 |  36 LGGC 151755    | 12/28/84  | C & P  | AJ   | N 3767268    SLOT 23
-------------------------------------------------------------------------------
  90 |  36 LGGS 90327     |  1/31/85  | C & P  | GS   | FDEA 379309  SLOT 24
-------------------------------------------------------------------------------
  91 |  359-2921          | 01/07/85  | C & P  |FRELIN| C 3771841 JAK 222
-------------------------------------------------------------------------------
  92 |  359-2922          | 01/07/85  | C & P  |FRELIN| C 3771841 JAK 223
-------------------------------------------------------------------------------
  93 |  359-2923          | 01/07/85  | C & P  |FRELIN| C 3771841 JAK 224
-------------------------------------------------------------------------------
  94 |  359-2924          | 01/07/85  | C & P  |FRELIN| C 3771841 JAK 227
-------------------------------------------------------------------------------
  95 |  359-2925          | 01/07/85  | C & P  |FRELIN| C 3771841 JAK 228
-------------------------------------------------------------------------------
  96 |  359-2926          | 01/07/85  | C & P  |FRELIN| C 3771841 JAK 229
-------------------------------------------------------------------------------
  97 |  359-2927          | 01/07/85  | C & P  |FRELIN| C 3771841 JAK 230
-------------------------------------------------------------------------------
  98 |  359-2928          | 01/07/85  | C & P  |FRELIN| C 3771841 JAK 231
-------------------------------------------------------------------------------
  99 |  359-2929          | 01/07/85  | C & P  |FRELIN| C 3771841 JAK 232
-------------------------------------------------------------------------------
 100 |  36 LGGS 151921    | 01/07/85  | C & P  | MTW  | FDEA 394523 SLOT 25
-------------------------------------------------------------------------------
 101 |  36 LGGC 154882    | 01/10/85  | C & P  | R    | N 3766884   SLOT 26
-------------------------------------------------------------------------------
 102 |  36 HCGS 81211 CV  | 01/10/85  | C & P  | R    | DHEA 339602 LL  T-1 BLOC
-------------------------------------------------------------------------------
 103 |  36 LGGC 155622    | 01/28/85  | C & P  | KRJ  | N 3770532    SLOT 27
-------------------------------------------------------------------------------
 104 |  36 LGGC 155623    | 01/28/85  | C & P  | KRJ  | C 3771387    SLOT 28
-------------------------------------------------------------------------------
 105 |  36 LGGC 155625    | 01/29/85  | C & P  | MTW  | N 3771390    SLOT 29
-------------------------------------------------------------------------------
 106 |                    |           |        |      |
-------------------------------------------------------------------------------
 107 |                    |           |        |      |
-------------------------------------------------------------------------------
 108 |                    |           |        |      |
-------------------------------------------------------------------------------
 109 |                    |           |        |      |
-------------------------------------------------------------------------------
 110 |                    |           |        |      |
-------------------------------------------------------------------------------
 